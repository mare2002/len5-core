// Copyright 2019 Politecnico di Torino.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 2.0 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-2.0. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// File: issue_decoder.sv
// Author: Michele Caon, Flavia Guella
// Date: 13/11/2019

module issue_decoder (
  // Instruction from the issue logic
  input len5_pkg::instr_t   instruction_i,  // the issuing instruction
  input csr_pkg::csr_priv_t priv_mode_i,    // current privilege mode

  // Issue decoder <--> issue CU
  output expipe_pkg::issue_type_t issue_type_o,  // issue operation type

  // Information to the issue logic
  output len5_pkg::except_code_t except_code_o,  // exception code to send to the ROB
  output expipe_pkg::issue_eu_t assigned_eu_o,  // assigned EU
  output logic skip_eu_o,  // do not assign to any EU
  output expipe_pkg::eu_ctl_t eu_ctl_o,  // controls for the assigned EU
  output logic mem_crit_o,  // memory accesses shall wait for this instruction to complete
  output logic order_crit_o,  // out-of-order commit not allowed
  output expipe_pkg::rs1_sel_t rs1_sel_o,  // rs1 source
  output expipe_pkg::rs2_sel_t rs2_sel_o,  // rs2 source
  output expipe_pkg::rs3_sel_t rs3_sel_o,  // rs3 source
  output logic rd_upd_o,  // the instruction updates a destination register rd
  output expipe_pkg::imm_format_t imm_format_o  // immediate format
);

  import len5_config_pkg::*;
  import len5_pkg::*;
  import expipe_pkg::*;
  import memory_pkg::*;
  import csr_pkg::*;
  import instr_pkg::*;

  // Parameters
  localparam logic [ILEN-1:0] RET = {12'b0, 5'b00001, 3'b000, 5'b00000, JALR[OPCODE_LEN-1:0]};

  // INTERNAL SIGNALS
  // ----------------
  // Exceptions
  except_code_t except_code;

  // Main decoder (opcode and special cases)
  issue_type_t  issue_type;
  issue_eu_t    assigned_eu;
  eu_ctl_t      eu_ctl;
  logic         mem_crit;  // stores must wait for these instruction completion
  logic         order_crit;  // out-of-order commit not allowed
  rs1_sel_t     rs1_sel;
  rs2_sel_t     rs2_sel;
  rs3_sel_t     rs3_sel;
  logic         rd_upd;
  imm_format_t  imm_format;
  logic         skip_eu;
  logic         opcode_except;

  // -------------------
  // INSTRUCTION DECODER
  // -------------------
  // New supported instructions can be added here. Instruction definitions
  // are taken from 'instr_pkg.sv', which is generated by the RISC-V opcode
  // generator called by 'sw/opcodes/gen_opcodes.sh'.

  // Main instruction decoder
  // ------------------------
  always_comb begin : main_decoder
    // Default values
    issue_type    = ISSUE_TYPE_NONE;
    skip_eu       = 1'b0;
    assigned_eu   = EU_INT_ALU;
    eu_ctl.raw    = '0;
    mem_crit      = 1'b1;  // opt-out policy is safer
    order_crit    = 1'b0;
    rs1_sel       = RS1_SEL_NONE;
    rs2_sel       = RS2_SEL_NONE;
    rs3_sel       = RS3_SEL_NONE;
    rd_upd        = 1'b1;  // true by default
    imm_format    = IMM_TYPE_I;
    opcode_except = 1'b0;
    except_code   = E_ILLEGAL_INSTRUCTION;

    // Main decoding logic
    unique casez (instruction_i.raw)
      // RV64I
      ADD: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_ADD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      ADDW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_ADDW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      ADDI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_ADD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      ADDIW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_ADDW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SUB: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SUB;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SUBW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SUBW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      AND: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_AND;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      ANDI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_AND;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      OR: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_OR;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      ORI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_OR;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      XOR: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_XOR;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      XORI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_XOR;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SLL: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLL;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SLLW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLLW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SLLI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLL;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SLLIW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLLW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SRL: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRL;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SRLW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRLW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SRLI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRL;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SRLIW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRLW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SRA: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRA;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SRAW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRAW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SRAI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRA;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SRAIW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SRAW;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SLT: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLT;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SLTU: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLTU;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
      end
      SLTI: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLT;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      SLTIU: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_SLTU;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_IMM;
      end
      LUI: begin
        issue_type = ISSUE_TYPE_LUI;
        skip_eu    = 1'b1;
        mem_crit   = 1'b0;
        imm_format = IMM_TYPE_U;
      end
      AUIPC: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_INT_ALU;
        eu_ctl.alu  = ALU_ADD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_PC;
        rs2_sel     = RS2_SEL_IMM;
        imm_format  = IMM_TYPE_U;
      end
      JAL: begin
        issue_type  = ISSUE_TYPE_JUMP;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = (instruction_i.j.rd == 5'b00001) ? BU_CALL : BU_JAL;
        mem_crit    = 1'b0;
        imm_format  = IMM_TYPE_J;
      end
      JALR: begin
        issue_type  = ISSUE_TYPE_JUMP;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = (instruction_i.raw == RET) ? BU_RET : BU_JALR;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      BEQ: begin
        issue_type  = ISSUE_TYPE_BRANCH;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = BU_BEQ;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_B;
      end
      BNE: begin
        issue_type  = ISSUE_TYPE_BRANCH;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = BU_BNE;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_B;
      end
      BLT: begin
        issue_type  = ISSUE_TYPE_BRANCH;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = BU_BLT;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_B;
      end
      BLTU: begin
        issue_type  = ISSUE_TYPE_BRANCH;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = BU_BLTU;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_B;
      end
      BGE: begin
        issue_type  = ISSUE_TYPE_BRANCH;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = BU_BGE;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_B;
      end
      BGEU: begin
        issue_type  = ISSUE_TYPE_BRANCH;
        assigned_eu = EU_BRANCH_UNIT;
        eu_ctl.bu   = BU_BGEU;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_B;
      end
      LB: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_BYTE;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      LBU: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_BYTE_U;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      LH: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_HALFWORD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      LHU: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_HALFWORD_U;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      LW: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_WORD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      LWU: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_WORD_U;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      LD: begin
        issue_type  = ISSUE_TYPE_INT;
        assigned_eu = EU_LOAD_BUFFER;
        eu_ctl.lsu  = LS_DOUBLEWORD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        imm_format  = IMM_TYPE_I;
      end
      SB: begin
        issue_type  = ISSUE_TYPE_STORE;
        assigned_eu = EU_STORE_BUFFER;
        eu_ctl.lsu  = LS_BYTE;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_S;
      end
      SH: begin
        issue_type  = ISSUE_TYPE_STORE;
        assigned_eu = EU_STORE_BUFFER;
        eu_ctl.lsu  = LS_HALFWORD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_S;
      end
      SW: begin
        issue_type  = ISSUE_TYPE_STORE;
        assigned_eu = EU_STORE_BUFFER;
        eu_ctl.lsu  = LS_WORD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_S;
      end
      SD: begin
        issue_type  = ISSUE_TYPE_STORE;
        assigned_eu = EU_STORE_BUFFER;
        eu_ctl.lsu  = LS_DOUBLEWORD;
        mem_crit    = 1'b0;
        rs1_sel     = RS1_SEL_INT;
        rs2_sel     = RS2_SEL_INT;
        rd_upd      = 1'b0;
        imm_format  = IMM_TYPE_S;
      end
      FENCE: begin
        issue_type = ISSUE_TYPE_STALL;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
      end
      ECALL: begin  // TODO: add ECALL support
        issue_type    = ISSUE_TYPE_EXCEPT;
        skip_eu       = 1'b1;
        order_crit    = 1'b1;
        opcode_except = 1'b1;
        unique case (priv_mode_i)
          PRIV_MODE_U: except_code = E_ENV_CALL_UMODE;
          PRIV_MODE_S: except_code = E_ENV_CALL_SMODE;
          default:     except_code = E_ENV_CALL_MMODE;
        endcase
      end
      EBREAK: begin  // TODO: add EBREAK support
        issue_type    = ISSUE_TYPE_EXCEPT;
        skip_eu       = 1'b1;
        order_crit    = 1'b1;
        opcode_except = 1'b1;
        except_code   = E_BREAKPOINT;
      end

      // RV64M
      MUL: begin
        if (LEN5_M_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_MULT;
          eu_ctl.mult = MULT_MUL;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      MULH: begin
        if (LEN5_M_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_MULT;
          eu_ctl.mult = MULT_MULH;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      MULHU: begin
        if (LEN5_M_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_MULT;
          eu_ctl.mult = MULT_MULHU;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      MULHSU: begin
        if (LEN5_M_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_MULT;
          eu_ctl.mult = MULT_MULHSU;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      MULW: begin
        if (LEN5_M_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_MULT;
          eu_ctl.mult = MULT_MULW;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      DIV: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_DIV;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      DIVU: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_DIVU;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      DIVW: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_DIVW;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      DIVUW: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_DIVUW;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      REM: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_REM;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      REMU: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_REMU;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      REMW: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_REMW;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      REMUW: begin
        if (LEN5_DIV_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_INT_DIV;
          eu_ctl.div  = DIV_REMUW;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end

      // RV32ZICSR
      // TODO: check CSR instructions
      CSRRW: begin
        issue_type = ISSUE_TYPE_CSR;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
        rs2_sel    = RS2_SEL_INT;
      end
      CSRRWI: begin
        issue_type = ISSUE_TYPE_CSR;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
        rs2_sel    = RS2_SEL_IMM;
      end
      CSRRS: begin
        issue_type = ISSUE_TYPE_CSR;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
        rs2_sel    = RS2_SEL_INT;
      end
      CSRRSI: begin
        issue_type = ISSUE_TYPE_CSR;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
        rs2_sel    = RS2_SEL_IMM;
      end
      CSRRC: begin
        issue_type = ISSUE_TYPE_CSR;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
        rs2_sel    = RS2_SEL_INT;
      end
      CSRRCI: begin
        issue_type = ISSUE_TYPE_CSR;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
        rs2_sel    = RS2_SEL_IMM;
      end

      // RV32SYSTEM
      // TODO: add support for SYSTEM instructions
      MRET: begin
        issue_type    = ISSUE_TYPE_EXCEPT;
        skip_eu       = 1'b1;
        order_crit    = 1'b1;
        opcode_except = 1'b1;
        except_code   = E_ENV_CALL_MMODE;
      end
      WFI: begin
        issue_type = ISSUE_TYPE_STALL;
        skip_eu    = 1'b1;
        order_crit = 1'b1;
      end

      // RV64F
      FLW: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_LOAD_BUFFER;
          eu_ctl.lsu  = LS_WORD;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          imm_format  = IMM_TYPE_I;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSW: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_STORE;
          assigned_eu = EU_STORE_BUFFER;
          eu_ctl.lsu  = LS_WORD;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_FP;
          rd_upd      = 1'b0;
          imm_format  = IMM_TYPE_S;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMADD_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MADD_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMSUB_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MSUB_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FNMSUB_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_NMSUB_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FNMADD_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_NMADD_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FADD_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_ADD_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSUB_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SUB_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMUL_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MUL_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FDIV_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_DIV_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSQRT_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SQRT_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSGNJ_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SGNJ_S;  // TODO: check, the actual op is distinguished through rm
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSGNJN_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SGNJ_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSGNJX_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SGNJ_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMIN_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MINMAX_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMAX_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MINMAX_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_W_S: begin  // single to int
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_S2I;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_WU_S: begin  // single to unsigned int
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_S2I_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_S_W: begin  // int to single
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_I2S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_S_WU: begin  // unsigned int to single
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_I2S_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_L_S: begin  // single to long int
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_S2L;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_LU_S: begin  // single to unsigned int
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_S2L_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_S_L: begin  // long to single
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_L2S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_S_LU: begin  // unsigned long to single
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_L2S_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMV_X_W: begin  // single to int
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_S2I;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMV_W_X: begin  // int to single
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_I2S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FEQ_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CMP_S;  // TODO: check, rm encodes comp type
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FLT_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CMP_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FLE_S: begin
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CMP_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCLASS_S: begin  // write to int RF
        if (LEN5_F_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CLASS_S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end

      // RV64D
      FLD: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_LOAD_BUFFER;
          eu_ctl.lsu  = LS_DOUBLEWORD;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          imm_format  = IMM_TYPE_I;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSD: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_STORE;
          assigned_eu = EU_STORE_BUFFER;
          eu_ctl.lsu  = LS_DOUBLEWORD;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_FP;
          rd_upd      = 1'b0;
          imm_format  = IMM_TYPE_S;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMADD_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MADD_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMSUB_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MSUB_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FNMSUB_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_NMSUB_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FNMADD_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_NMADD_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
          rs3_sel     = RS3_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FADD_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_ADD_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSUB_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SUB_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMUL_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MUL_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FDIV_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_DIV_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSQRT_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SQRT_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSGNJ_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SGNJ_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSGNJN_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SGNJ_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FSGNJX_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_SGNJ_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMIN_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MINMAX_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMAX_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_MINMAX_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_S_D: begin  // double to single
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_D2S;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_D_S: begin  // single to double
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_S2D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_W_D: begin  // double to int
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_D2I;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_WU_D: begin  // double to 32-bit int
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_D2I_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_D_W: begin  //32-bit int to double
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_I2D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_D_WU: begin  // unsigned 32-bit int to double
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_I2D_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_L_D: begin  // double to 64-bit int
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_D2L;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_LU_D: begin  // double to 64-bit unsigned int
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_D2L_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_D_L: begin  // long int to double
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_L2D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCVT_D_LU: begin  // unsigned long int to double
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_L2D_U;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMV_X_D: begin  // double to 64-bit int
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_D2L;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FMV_D_X: begin  // int to fp reg
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_FP;  // FP RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_L2D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FEQ_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CMP_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FLT_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CMP_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FLE_D: begin
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CMP_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
          rs2_sel     = RS2_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      FCLASS_D: begin  // write to int RF
        if (LEN5_D_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_FPU;
          eu_ctl.fpu  = FPU_CLASS_D;  // TODO: check
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_FP;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end

      // DUMMY COPR
      XDUMMY_ITERATIVE: begin
        if (LEN5_DUMMY_COPR_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;  // int RF destination
          assigned_eu = EU_DUMMY_COPR;
          eu_ctl.copr = DUMMY_ITERATIVE;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_IMM;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      XDUMMY_PIPE: begin
        if (LEN5_DUMMY_COPR_EN != 1'b0) begin
          issue_type  = ISSUE_TYPE_INT;
          assigned_eu = EU_DUMMY_COPR;
          eu_ctl.copr = DUMMY_PIPELINE;
          mem_crit    = 1'b0;
          rs1_sel     = RS1_SEL_INT;
          rs2_sel     = RS2_SEL_IMM;
        end else begin
          issue_type    = ISSUE_TYPE_EXCEPT;
          skip_eu       = 1'b1;
          opcode_except = 1'b1;
        end
      end
      // Unsupported instruction
      default: begin
        issue_type    = ISSUE_TYPE_EXCEPT;
        skip_eu       = 1'b1;
        opcode_except = 1'b1;
      end
    endcase
  end

  assign issue_type_o  = (opcode_except) ? ISSUE_TYPE_EXCEPT : issue_type;
  assign skip_eu_o     = (opcode_except) ? 1'b1 : skip_eu;

  // -----------------
  // OUTPUT GENERATION
  // -----------------
  assign except_code_o = except_code;
  assign assigned_eu_o = assigned_eu;
  assign eu_ctl_o      = eu_ctl;
  assign mem_crit_o    = mem_crit;
  assign order_crit_o  = order_crit;
  assign rs1_sel_o     = rs1_sel;
  assign rs2_sel_o     = rs2_sel;
  assign rs3_sel_o     = rs3_sel;
  assign rd_upd_o      = rd_upd;
  assign imm_format_o  = imm_format;

  // ----------
  // ASSERTIONS
  // ----------
`ifndef SYNTHESIS
`ifndef VERILATOR
  /* Assertions here */
`endif  /* VERILATOR */
`endif  /* SYNTHESIS */

endmodule
